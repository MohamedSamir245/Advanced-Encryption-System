function [31:0] RotWord_fn(input [31:0]word);


RotWord_fn={word[23:0],word[31:24]};
endfunction
